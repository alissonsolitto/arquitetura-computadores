LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY RAM IS
    PORT ( CLK  : IN  STD_LOGIC;
           RST  : IN  STD_LOGIC;
		   ADDR : IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
           RW   : IN  STD_LOGIC;
           DIN  : IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
           DOUT : OUT  STD_LOGIC_VECTOR (7 DOWNTO 0));
END RAM;

ARCHITECTURE BEHAVIORAL OF RAM IS
TYPE RAM_TYPE IS ARRAY(0 TO 255) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL RAM: RAM_TYPE;

BEGIN
   PROCESS(CLK, RST) IS
	BEGIN
	   IF (RST = '1') THEN

			RAM(0) <= "10100001"; -- A1 - LE O NUMERO 1
			RAM(1) <= "10100010"; -- A2 - LE O NUMERO 2
			RAM(2) <= "10100011"; -- A3 - LE O OPERADOR			
			RAM(3) <= "10111011"; -- BB - EFETUA A OPERACAO
			RAM(4) <= "11001100"; -- CC - MOSTRA VALOR NO DISPLAY
			
					
		ELSIF CLK'EVENT AND CLK = '1' THEN
			IF(RW = '1') THEN -- ESCREVER NA MEMORIA
			  RAM(TO_INTEGER(UNSIGNED(ADDR))) <= DIN;			
			END IF;			
		END IF;
		
	END PROCESS;
	
	-- N�O PRECISA DE CLOCK PARA LER NA MEMORIA
	DOUT <= RAM(TO_INTEGER(UNSIGNED(ADDR)));
	
END BEHAVIORAL;
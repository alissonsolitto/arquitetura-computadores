LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY PISCA IS
    PORT ( CLK : IN  STD_LOGIC;
           LED : OUT  STD_LOGIC);
END PISCA;

ARCHITECTURE BEHAVIORAL OF PISCA IS
SIGNAL CONT: INTEGER RANGE 0 TO 300000001;
BEGIN
  PROCESS (CLK)
  BEGIN
    IF CLK'EVENT AND CLK='1' THEN
	   
		CONT <= CONT + 1;
		
		IF(CONT <=  200000000) THEN
		  LED <= '0';
		ELSE
        LED <= '1';
		END IF;
		
		IF CONT = 300000000 THEN
		  CONT <=0;
		END IF;
	 
	 END IF;
	 
  END PROCESS;


END BEHAVIORAL;
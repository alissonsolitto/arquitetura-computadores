LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TOP IS
    PORT ( CLK : IN  STD_LOGIC;
           RST : IN  STD_LOGIC;			     
           ENTER: IN STD_LOGIC;
  	        OPER : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
           NUM  : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			  AN   : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			  SEG  : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);			  
           LED : OUT  STD_LOGIC_VECTOR (7 DOWNTO 0));
END TOP;

ARCHITECTURE BEHAVIORAL OF TOP IS
--COMPONENTE RAM
COMPONENT RAM IS
    PORT ( CLK  : IN  STD_LOGIC;
           RST  : IN  STD_LOGIC;
           ADDR : IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
           RW   : IN  STD_LOGIC;
           DIN  : IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
           DOUT : OUT  STD_LOGIC_VECTOR (7 DOWNTO 0));
END COMPONENT;

--COMPONENTE HC05
COMPONENT HC05 IS
    PORT ( 	CLK  : IN  STD_LOGIC;
			RST  : IN  STD_LOGIC;
			ENTER: IN STD_LOGIC;
			OPER : IN STD_LOGIC_VECTOR (1 DOWNTO 0);			  
			NUM  : IN STD_LOGIC_VECTOR (3 DOWNTO 0);				   
			DOUT : IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
			ADDR : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			RW   : OUT STD_LOGIC;
			DIN  : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);			  
			AN   : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			SEG  : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
			LED  : OUT  STD_LOGIC_VECTOR (7 DOWNTO 0));
END COMPONENT;

--SINAIS
SIGNAL DOUT : STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL ADDR : STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL RW   : STD_LOGIC;
SIGNAL DIN  : STD_LOGIC_VECTOR (7 DOWNTO 0);

SIGNAL CONT: INTEGER RANGE 0 TO 100000001; -- 1S
SIGNAL CLOCK_DIV: STD_LOGIC;

BEGIN
  --MAPEANDO COMPONENTES
  RAM1 : RAM  PORT MAP(CLOCK_DIV, RST, ADDR, RW, DIN, DOUT);
  HC051: HC05 PORT MAP(CLOCK_DIV, RST, ENTER, OPER, NUM, DOUT, ADDR, RW, DIN, AN, SEG, LED);
  
   PROCESS(CLK, RST) IS
	BEGIN
	   IF (RST = '1') THEN
			CONT <= 0;
		ELSIF CLK'EVENT AND CLK = '1' THEN		
			CONT <= CONT + 1;
			IF(CONT <= 500000)THEN
				CLOCK_DIV <= '0';
			ELSE	
				CLOCK_DIV <= '1';
			END IF;	
			
			IF(CONT = 1000000)THEN
				CONT <= 0;
			END IF;
		END IF;
	END PROCESS;  


END BEHAVIORAL;